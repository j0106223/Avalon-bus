module clk_gen (
    clk_i,
    clk_o
);
    input clk_i;
    output clk_o;
    
endmodule