`default_nettype none
module i2c_core (
    clk,
    reset_n,
    sda,
    scl,
);
    input clk;
    input reset_n; 
endmodule