module dma_core (
    clk,
    reset_n,
    data_i,
    data_o,
);
    localparam IDLE;
    localparam DONE;
//=============FSM===============
//=============FSM===============
endmodule