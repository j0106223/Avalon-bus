module rv32_single (
    address,
    data,
);
    //instruction master
    //data master
endmodule