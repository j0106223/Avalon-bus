`default_nettype none
module rv32_5stage (
    address,
    data,

);
    output address;
    //instruction master
    //data master
endmodule