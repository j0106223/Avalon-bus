module x_dec (
    ports
);
    
endmodule