module ps2_core (
    clk,
    reset_n,
    sclk,
    data
);
    
endmodule