module i2s_core (
    clk,
    reset_n,
);
    input clk;
    input reset_n;    
endmodule