module avs_i2s (
    clk,
    reset_n,
    avs_s0_address,
    avs_s0_read,
    avs_s0_write,
    avs_s0_waitrequest,
    avs_s0_readdata,
    avs_s0_writedata
);
    input clk;
    input reset_n;
    input        avs_s0_address;
    input        avs_s0_read;
    input        avs_s0_write;
    output       avs_s0_waitrequest;
    output [31:0]avs_s0_readdata;
    input  [31:0]avs_s0_writedata;

//==================register map begin======================

//==================register map end========================
    //write register
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)begin

        end else begin
            if(avs_s0_write)begin
                case (avs_s0_address)
                    0:
                    0:
                    0:
                    0: 
                    default:begin
                    end 
                endcase
            end
        end
    end

    always @(*) begin
        if(avs_s0_read)begin
            case (avs_s0_address)
                : 
                default:begin
                end
            endcase
        end
    end

    wire i2s_clk;

    i2s_core i2s_core_inst(
        .reset_n(reset_n),
        .data_right(),
        .data_left(),
        .sck(i2s_clk),
        .sd(),
        .ws()
    );

    clk_gen clk_gen_i2s(
        .clk_i   (clk),
        .reset_n (reset_n),
        .clk_div (clk_div),
        .clk_o   (i2s_clk)
    );
endmodule