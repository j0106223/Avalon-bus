module avs_uare_tb;
    


    
endmodule