module top (

);
    
endmodule