module sim_top (
    clk,
    reset_n,
    sim_clk,
    sim_reset_n,
    sim_io
);

    input  clk;
    input  reset_n;
    output sim_clk;
    output sim_reset_n;
    inout  sim_io;

      
endmodule